module fruit_check(
	input [9:0] x0,		//Centre of Fruit
	input [9:0] y0,		//Centre of Fruit
	input [9:0] x,		//Co-ordinate to be tested
	input [9:0] y,		//Co-ordinate to be tested
	input [1:0] choice,	//Fruit choice
	input en,			//ENABLE
	input clk,			//CLOCK
	output [11:0] color	//Color to display
	
);

	reg [9:0] xt;
	reg [9:0] yt;
	reg [9:0] int_x;
	reg [9:0] int_y;
	reg [11:0] fruit_color;
 	reg ch;

	assign int_x = x0 >> 0;
	assign int_y = y0 >> 0;	

	assign xt = (x > int_x) ? x - int_x : int_x - x ;

	always @ (posedge clk)
	begin

	assign yt = y - int_y + 10'b0000001000 ;
	
	case (choice)

	2'b00:	//ORANGE
		begin 
		assign fruit_color = 12'b111110001000 ;
		
		case (yt) 
			10'b0000000000 : ch = (xt < 10'b0000000011) ? 1'b1 : 1'b0 ; 
			10'b0000000001 : ch = (xt < 10'b0000000101) ? 1'b1 : 1'b0 ;
			10'b0000000010 : ch = (xt < 10'b0000000110) ? 1'b1 : 1'b0 ;
			10'b0000000011 : ch = (xt < 10'b0000000111) ? 1'b1 : 1'b0 ;
			10'b0000000100 : ch = (xt < 10'b0000001000) ? 1'b1 : 1'b0 ;
			10'b0000000101 : ch = (xt < 10'b0000001000) ? 1'b1 : 1'b0 ;
			10'b0000000110 : ch = (xt < 10'b0000001001) ? 1'b1 : 1'b0 ;
			10'b0000000111 : ch = (xt < 10'b0000001001) ? 1'b1 : 1'b0 ;
			10'b0000001000 : ch = (xt < 10'b0000001001) ? 1'b1 : 1'b0 ;
			10'b0000001001 : ch = (xt < 10'b0000001001) ? 1'b1 : 1'b0 ;
			10'b0000001010 : ch = (xt < 10'b0000001001) ? 1'b1 : 1'b0 ;
			10'b0000001011 : ch = (xt < 10'b0000001000) ? 1'b1 : 1'b0 ;
			10'b0000001100 : ch = (xt < 10'b0000001000) ? 1'b1 : 1'b0 ;
			10'b0000001101 : ch = (xt < 10'b0000000111) ? 1'b1 : 1'b0 ;
			10'b0000001110 : ch = (xt < 10'b0000000110) ? 1'b1 : 1'b0 ;
			10'b0000001111 : ch = (xt < 10'b0000000101) ? 1'b1 : 1'b0 ;
			10'b0000010000 : ch = (xt < 10'b0000000011) ? 1'b1 : 1'b0 ;
		endcase
		end

	2'b01:	//APPLE
		begin 
		assign fruit_color = 12'b111100000000 ;
	
		case (yt) 
			10'b0000000000 : ch = (xt < 10'b0000000001) ? 1'b1 : 1'b0 ;
			10'b0000000001 : ch = ((xt > 10'b0000000001 && xt < 10'b0000000111) || xt < 10'b0000000001) ? 1'b1 : 1'b0 ;
			10'b0000000010 : ch = (xt < 10'b0000001000) ? 1'b1 : 1'b0 ;
			10'b0000000011 : ch = (xt < 10'b0000001001) ? 1'b1 : 1'b0 ;
			10'b0000000100 : ch = (xt < 10'b0000001001) ? 1'b1 : 1'b0 ;
			10'b0000000101 : ch = (xt < 10'b0000001001) ? 1'b1 : 1'b0 ;
			10'b0000000110 : ch = (xt < 10'b0000001001) ? 1'b1 : 1'b0 ;
			10'b0000000111 : ch = (xt < 10'b0000001001) ? 1'b1 : 1'b0 ;
			10'b0000001000 : ch = (xt < 10'b0000001001) ? 1'b1 : 1'b0 ;
			10'b0000001001 : ch = (xt < 10'b0000001001) ? 1'b1 : 1'b0 ; 
			10'b0000001010 : ch = (xt < 10'b0000001001) ? 1'b1 : 1'b0 ; 
			10'b0000001011 : ch = (xt < 10'b0000001001) ? 1'b1 : 1'b0 ; 
			10'b0000001100 : ch = (xt < 10'b0000001001) ? 1'b1 : 1'b0 ; 
			10'b0000001101 : ch = (xt < 10'b0000001000) ? 1'b1 : 1'b0 ; 
			10'b0000001110 : ch = (xt < 10'b0000001000) ? 1'b1 : 1'b0 ; 
			10'b0000001111 : ch = (xt > 10'b0000000001 && xt < 10'b0000000111) ? 1'b1 : 1'b0 ; 
			10'b0000010000 : ch = (xt > 10'b0000000011 && xt < 10'b0000000110) ? 1'b1 : 1'b0 ; 
		endcase
		end
	
	2'b10:	//POMEGRANATE
		begin 
		assign fruit_color = 12'b111110111110 ;

		case (yt) 
			10'b0000000000 : ch = (xt == 10'b0000000011) ? 1'b1 : 1'b0 ;
			10'b0000000001 : ch = (xt > 10'b0000000000 && xt < 10'b0000000011) ? 1'b1 : 1'b0 ;
			10'b0000000010 : ch = (xt < 10'b0000000101) ? 1'b1 : 1'b0 ;
			10'b0000000011 : ch = (xt < 10'b0000000111) ? 1'b1 : 1'b0 ;
			10'b0000000100 : ch = (xt < 10'b0000001000) ? 1'b1 : 1'b0 ;
			10'b0000000101 : ch = (xt < 10'b0000001001) ? 1'b1 : 1'b0 ;
			10'b0000000110 : ch = (xt < 10'b0000001001) ? 1'b1 : 1'b0 ;
			10'b0000000111 : ch = (xt < 10'b0000001001) ? 1'b1 : 1'b0 ;
			10'b0000001000 : ch = (xt < 10'b0000001001) ? 1'b1 : 1'b0 ;
			10'b0000001001 : ch = (xt < 10'b0000001001) ? 1'b1 : 1'b0 ;
			10'b0000001010 : ch = (xt < 10'b0000001001) ? 1'b1 : 1'b0 ; 
			10'b0000001011 : ch = (xt < 10'b0000001001) ? 1'b1 : 1'b0 ; 
			10'b0000001100 : ch = (xt < 10'b0000001000) ? 1'b1 : 1'b0 ; 
			10'b0000001101 : ch = (xt < 10'b0000000111) ? 1'b1 : 1'b0 ; 
			10'b0000001110 : ch = (xt < 10'b0000000110) ? 1'b1 : 1'b0 ; 
			10'b0000001111 : ch = (xt < 10'b0000000101) ? 1'b1 : 1'b0 ; 
			10'b0000010000 : ch = (xt < 10'b0000000011) ? 1'b1 : 1'b0 ; 
		endcase
		end

	2'b11:	//PEAR
		begin 
		assign fruit_color = 12'b100111110000 ;

		case (yt) 
			10'b0000000000 : ch = (xt < 10'b0000000010) ? 1'b1 : 1'b0 ;
			10'b0000000001 : ch = (xt < 10'b0000000011) ? 1'b1 : 1'b0 ;
			10'b0000000010 : ch = (xt < 10'b0000000011) ? 1'b1 : 1'b0 ;
			10'b0000000011 : ch = (xt < 10'b0000000100) ? 1'b1 : 1'b0 ;
			10'b0000000100 : ch = (xt < 10'b0000000100) ? 1'b1 : 1'b0 ;
			10'b0000000101 : ch = (xt < 10'b0000000100) ? 1'b1 : 1'b0 ;
			10'b0000000110 : ch = (xt < 10'b0000000100) ? 1'b1 : 1'b0 ;
			10'b0000000111 : ch = (xt < 10'b0000000101) ? 1'b1 : 1'b0 ;
			10'b0000001000 : ch = (xt < 10'b0000000101) ? 1'b1 : 1'b0 ;
			10'b0000001001 : ch = (xt < 10'b0000000110) ? 1'b1 : 1'b0 ; 
			10'b0000001010 : ch = (xt < 10'b0000000111) ? 1'b1 : 1'b0 ; 
			10'b0000001011 : ch = (xt < 10'b0000000111) ? 1'b1 : 1'b0 ; 
			10'b0000001100 : ch = (xt < 10'b0000000111) ? 1'b1 : 1'b0 ; 
			10'b0000001101 : ch = (xt < 10'b0000000111) ? 1'b1 : 1'b0 ; 
			10'b0000001110 : ch = (xt < 10'b0000000111) ? 1'b1 : 1'b0 ; 
			10'b0000001111 : ch = (xt < 10'b0000000110) ? 1'b1 : 1'b0 ; 
			10'b0000010000 : ch = (xt < 10'b0000000100) ? 1'b1 : 1'b0 ; 
		endcase
		end

	assign color = (ch & en) ? fruit_color : 12'b0 ; 

	endcase
	
	end   
		
endmodule // FRUIT_CHECK
